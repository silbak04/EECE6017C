library verilog;
use verilog.vl_types.all;
entity shift_reg_tb is
end shift_reg_tb;
