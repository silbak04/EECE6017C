/*--==========================================================================--*/
//--================================ VERILOG ===================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: shift_register.v                                                --
//--                                                                            --
//-- DATE: 9/10/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: 4 bit shift register                                          --
//--                                                                            --
//--============================================================================--
//--================================ VERILOG ===================================--
/*--===========================================================================--*/

module shift_register (
    input clk, rst, d,
    output reg [3:0] shift_reg = 4'b0000
);

    always @ (posedge clk) begin
        if(rst)
            shift_reg <= 4'b0000;
        else
            shift_reg [3:1] <= shift_reg [2:0];
            shift_reg [0] <= d;
    end

endmodule
