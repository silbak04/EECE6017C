/*--==========================================================================--*/
//--================================ VERILOG ===================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: top.v                                                       --
//--                                                                            --
//-- DATE: 9/10/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: top module to instantiate flip flop and d latch               --
//--                                                                            --
//--============================================================================--
//--================================ VERILOG ===================================--
/*--===========================================================================--*/

module top (
    input clk, d,
    output q_a, q_b, q_c
);

    d_latch gated (
        .clk(clk),
        .d(d),
        .q_out(q_a)
    );

    flip_flop positive (
        .clk(clk),
        .d(d),
        .q_out(q_b)
    );

    flip_flop negative (
        .clk(~clk),
        .d(d),
        .q_out(q_c)
    );

endmodule
