/*--==========================================================================--*/
//--================================ VERILOG ===================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: d_latch.v                                                       --
//--                                                                            --
//-- DATE: 9/10/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: d latch                                                       --
//--                                                                            --
//--============================================================================--
//--================================ VERILOG ===================================--
/*--===========================================================================--*/

module d_latch (
    input clk, d,
    output q_out
);

    wire R_g, S_g, q, q_not; /* synthesis keep */ 

    nand (R_g, ~d, clk);
    nand (S_g, d, clk);
    nand (q, q_not, S_g);
    nand (q_not, q, R_g);

    assign q_out = q;

endmodule
