library verilog;
use verilog.vl_types.all;
entity rs_latch_tb is
end rs_latch_tb;
