library verilog;
use verilog.vl_types.all;
entity fsm_tb is
end fsm_tb;
