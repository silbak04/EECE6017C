/*--==========================================================================--*/
//--================================= VERILOG ==================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: d_fflop.v                                                       --
//--                                                                            --
//-- DATE: 9/10/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: d flip flop                                                   --
//--                                                                            --
//--============================================================================--
//--================================= VERILOG ==================================--
/*--===========================================================================--*/

module d_fflop (
    input clk, rst, d,
    output reg q_out = 0
);
    
    always @ (posedge clk) begin
        if(rst)
            q_out <= 0;
        else
            q_out <= d;
    end
endmodule
