library verilog;
use verilog.vl_types.all;
entity d_latch_tb is
end d_latch_tb;
