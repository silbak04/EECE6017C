/*--==========================================================================--*/
//--================================ VERILOG ===================================--
//--============================================================================--
//--                                                                            --
//-- FILE NAME: rs_latch.v                                                      --
//--                                                                            --
//-- DATE: 9/10/2012                                                            --
//--                                                                            --
//-- DESIGNER: Samir Silbak                                                     --
//--           silbak04@gmail.com                                               --
//--                                                                            --
//-- DESCRIPTION: rs latch                                                      --
//--                                                                            --
//--============================================================================--
//--================================ VERILOG ===================================--
/*--===========================================================================--*/

module rs_latch (
    input clk, R, S,
    output q_out
);

    wire R_g, S_g, q, q_not; /* synthesis keep */ 

    and (R_g, R, clk);
    and (S_g, S, clk);
    nor (q, R_g, q_not);
    nor (q_not, S_g, q);

    assign q_out = q;

endmodule
